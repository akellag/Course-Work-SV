module data(clk, reset, start, prod_reg_ld_high, prod_reg_shift_rt_a, prod_reg_shift_rt_b, )